--------------------------------------------------------------------------
-- Arquivo   : genius_musical_tb.vhd
-- Projeto   : Experiencia 06 - Projeto Base do Jogo do Desafio da Memória
--------------------------------------------------------------------------
-- Descricao : testbench para simulação com ModelSim
--
--             Cenário: Jogador vence
--             
--------------------------------------------------------------------------
-- Revisoes  :
--     Data        Versao  Autor             Descricao
--     01/02/2020  1.0     João Pedro C.M.   criacao
--------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

-- entidade do testbench
entity genius_musical_tb is
end entity;

architecture tb of genius_musical_tb is

  -- Componente a ser testado (Device Under Test -- DUT)
  component genius_musical is
    port (
      clock     : in  std_logic;
      reset     : in  std_logic;
      iniciar   : in  std_logic;
      ativar    : in  std_logic;
      botoes    : in  std_logic_vector(3 downto 0);
      notas     : out std_logic_vector(3 downto 0);
      jogador   : out std_logic;
      ganhou    : out std_logic;
      perdeu    : out std_logic;
      db_jogada                : out std_logic_vector(6 downto 0);
      db_rodada                : out std_logic_vector(6 downto 0);
      db_contagem              : out std_logic_vector(6 downto 0);
      db_memoria               : out std_logic_vector(6 downto 0);
      db_estado                : out std_logic_vector(6 downto 0)
    );
  end component;
  
  ---- Declaracao de sinais de entrada para conectar o componente
  signal clk_in     : std_logic := '0';
  signal rst_in     : std_logic := '0';
  signal iniciar_in : std_logic := '0';
  signal botoes_in  : std_logic_vector(3 downto 0) := "0000";
  signal ativar_in  : std_logic := '0';

  ---- Declaracao dos sinais de saida
  signal ganhou_out     : std_logic := '0';
  signal perdeu_out     : std_logic := '0';
  signal jogador_out    : std_logic := '0';
  signal notas_out      : std_logic_vector(3 downto 0);
  signal contagem_out   : std_logic_vector(6 downto 0) := "0000000";
  signal memoria_out    : std_logic_vector(6 downto 0);
  signal jogada_out     : std_logic_vector(6 downto 0);
  signal estado_out     : std_logic_vector(6 downto 0) := "0000000";
  signal rodada_out     : std_logic_vector(6 downto 0);

  -- Configurações do clock
  signal keep_simulating: std_logic := '0'; -- delimita o tempo de geração do clock
  constant clockPeriod : time := 20 ns;     -- frequencia 100MHz

  -- Configuração de jogo
  constant rodada : natural := 16; -- Nível de dificuldade
  constant modo   : natural := 3;

  -- Array de testes
  type   test_vector is array(0 to 15) of std_logic_vector(3 downto 0);
  signal tests : test_vector := (
                                   --C_Major ? (AINDA EM DEBATE)
                                   "0001", --G5 (783.99 Hz)
                                   "0010", --F5
                                   "0011", --E5
                                   "0100", --D5
                                   "0101", --C5 (523.25 Hz)
                                   "0110", --B5
                                   "0111", --A5
                                   "1000", --G4
                                   "1001", --F4
                                   "1010", --E4
                                   "1011", --D4
                                   "1100", --C4 (261.63 Hz) 
                                   "1011", --D4
                                   "1010", --E4
                                   "1001", --F4
                                   "1000");--G4
  
begin
  -- Gerador de clock: executa enquanto 'keep_simulating = 1', com o período especificado. 
  -- Quando keep_simulating=0, clock é interrompido, bem como a simulação de eventos
  clk_in <= (not clk_in) and keep_simulating after clockPeriod/2;
  
  ---- DUT para Simulacao
  DUT: genius_musical
       port map (
          clock           => clk_in,
          reset           => rst_in,
          iniciar         => iniciar_in,
          ativar          => ativar_in,
          botoes          => botoes_in,
          ganhou          => ganhou_out,
          perdeu          => perdeu_out,
          jogador         => jogador_out,
          notas           => notas_out,
          db_jogada       => jogada_out,
          db_contagem     => contagem_out,
          db_estado       => estado_out,
          db_memoria      => memoria_out,
          db_rodada       => rodada_out
       );
 
  ---- Gera sinais de estimulo para a simulacao
  stimulus: process is
  begin

    -- inicio da simulacao
    assert false report "inicio da simulacao" severity note;
    keep_simulating <= '1';  -- inicia geracao do sinal de clock

    ativar_in <= '0';
    -- gera pulso de reset (1 periodo de clock)
    rst_in <= '1';
    wait for clockPeriod;
    rst_in <= '0';

    -- espera para inicio dos testes
    wait for 10*clockPeriod;
    wait until falling_edge(clk_in);

    -- pulso do sinal de Iniciar (muda na borda de descida do clock)
    wait until falling_edge(clk_in);
    iniciar_in <= '1';
    wait until falling_edge(clk_in);
    iniciar_in <= '0';
    wait for 10*clockPeriod;
    -- Escolher Modo
    botoes_in  <= std_logic_vector(to_unsigned(modo, 4));
    ativar_in   <= '1';
    wait for 10*clockPeriod;
    botoes_in  <= "0000";
    ativar_in   <= '0'; 
    wait for 2*clockPeriod;
    -- Escolher Dificuldade
    botoes_in  <= std_logic_vector(to_unsigned(rodada-1, 4));
    ativar_in   <= '1';
    wait for 10*clockPeriod;
    ativar_in   <= '0'; 
    botoes_in  <= "0000";
    wait for 505*clockPeriod;
    tests(0) <= notas_out;
    assert ganhou_out   = '0'    report "bad initial ganhou"                      severity error;
    assert perdeu_out   = '0'    report "bad initial perdeu"                      severity error;
    wait for 500*clockPeriod;
    -- Cada iteração corresponde a uma rodada
    for i in 0 to rodada - 1 loop
      assert false report "Rodada " & integer'image(i) severity note;
      -- Cada iteração corresponde a uma jogada
      -- Última rodada -> sem escrita
      if(i = rodada - 1) then
        for k in 0 to i loop 
          botoes_in  <= tests(k);
          ativar_in   <= '1';
          wait for 3*clockPeriod;
          assert notas_out = tests(k) report "bad nota = " & integer'image(to_integer(unsigned(notas_out))) severity error;
          -- última jogada da última rodada -> ganhou!
            assert ganhou_out   = '0'  report "bad ganhou"                          severity error;
            assert perdeu_out   = '0'  report "bad perdeu"                          severity error;
            wait for 9*clockPeriod;
            botoes_in  <= "0000";
            ativar_in   <= '0';
            wait for 3*clockPeriod;
            assert notas_out     = "0000"   report "bad nota = " & integer'image(to_integer(unsigned(notas_out))) severity error;
            if(k = rodada - 1) then
              assert ganhou_out   = '1'  report "bad ganhou"  severity error;
              assert perdeu_out   = '0'  report "bad perdeu"  severity error;
            else
              assert ganhou_out   = '0' report "bad ganhou"   severity error;
              assert perdeu_out   = '0' report "bad perdeu"   severity error;
            end if;
            wait for 9*clockPeriod;
        end loop;
      -- Demais rodadas -> escrita pós-jogada
      else
        for k in 0 to i + 1 loop 
          if(k = i + 1) then
            -- Modo multijogador -> jogador escreve a próxima jogada
            if(modo = 2) then
              botoes_in  <= tests(k);
              ativar_in   <= '1';
              wait for 3*clockPeriod;
              assert notas_out     = tests(k) report "bad nota = " & integer'image(to_integer(unsigned(notas_out))) severity error;
            -- Demais modos -> jogador ve a jogada, determinada pela FPGA, e imita ela
            else
              wait for 500*clockPeriod;
              tests(k) <= notas_out;
              wait for 250*clockPeriod;
              assert notas_out     = tests(k) report "bad nota = " & integer'image(to_integer(unsigned(notas_out))) severity error;
              wait for 253*clockPeriod;
            end if;
          else
            botoes_in <= tests(k);
            ativar_in  <= '1';
            wait for 3*clockPeriod;
            assert notas_out     = tests(k) report "bad nota = " & integer'image(to_integer(unsigned(notas_out))) severity error;
          end if;
          assert ganhou_out   = '0'      report "bad  ganhou"                             severity error;
          assert perdeu_out   = '0'      report "bad  perdeu"                             severity error;
          wait for 9*clockPeriod;
          botoes_in  <= "0000";
          ativar_in   <= '0';
          wait for 3*clockPeriod;
          assert ganhou_out   = '0'      report "bad  ganhou"                             severity error;
          assert perdeu_out   = '0'      report "bad  perdeu"                             severity error;
          wait for 9*clockPeriod;
        end loop;
      end if;
    end loop;

    ---- final do testbench
    assert false report "fim da simulacao" severity note;
    keep_simulating <= '0';
    
    wait; -- fim da simulação: processo aguarda indefinidamente
  end process;

end architecture;